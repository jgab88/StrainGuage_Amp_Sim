** Profile: "SCHEMATIC1-StrainResponse"  [ d:\users\jerryg\projects\pspice_practice\first_ws\StrainGuage_Amp\StrainGuage_Amp-PSpiceFiles\SCHEMATIC1\StrainResponse.sim ] 

** Creating circuit file "StrainResponse.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM Rgauge 315 385 5 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ABSTOL= 1e-6
.OPTIONS ITL4= 50
.OPTIONS RELTOL= 0.01
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
