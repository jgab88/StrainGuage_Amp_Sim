** Profile: "SCHEMATIC1-Rgauge"  [ d:\users\jerryg\projects\pspice_practice\first_ws\StrainGuage_Amp\StrainGuage_Amp-PSpiceFiles\SCHEMATIC1\Rgauge.sim ] 

** Creating circuit file "Rgauge.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM Rgauge 350 360 1 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ITL4= 50
.OPTIONS THREADS= 36
.OPTIONS PTRANABSTOL= 1e-5
.OPTIONS PTRANVNTOL= 1e-4
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
